module BDC_7SEGx(
    input [27:0] code,
    input CLK,
    output reg [7:0] BCD0, BCD1, BCD2, BCD3, BCD4, BCD5, BCD6
);

initial begin
    BCD0 = 7'b0111111;
    BCD1 = 7'b0111111;
    BCD2 = 7'b0111111;
    BCD3 = 7'b0111111;
    BCD4 = 7'b0111111;
    BCD5 = 7'b0111111;
    BCD6 = 7'b0111111;
end

always @ (posedge CLK) begin
        case(code[3:0])
            4'b0000: BCD0 = 7'b1000000;
            4'b0001: BCD0 = 7'b1111001;
            4'b0010: BCD0 = 7'b0100100;
            4'b0011: BCD0 = 7'b0110000;
            4'b0100: BCD0 = 7'b0011001;
            4'b0101: BCD0 = 7'b0010010;
            4'b0110: BCD0 = 7'b0000010;
            4'b0111: BCD0 = 7'b1111000;
            4'b1000: BCD0 = 7'b0000000;
            4'b1001: BCD0 = 7'b0011000;
            4'b1010: BCD0 = 7'b0111111;
        endcase
        case(code[7:4])
            4'b0000: BCD1 = 7'b1000000;
            4'b0001: BCD1 = 7'b1111001;
            4'b0010: BCD1 = 7'b0100100;
            4'b0011: BCD1 = 7'b0110000;
            4'b0100: BCD1 = 7'b0011001;
            4'b0101: BCD1 = 7'b0010010;
            4'b0110: BCD1 = 7'b0000010;
            4'b0111: BCD1 = 7'b1111000;
            4'b1000: BCD1 = 7'b0000000;
            4'b1001: BCD1 = 7'b0011000;
            4'b1010: BCD1 = 7'b0111111;
        endcase
        case(code[11:8])
            4'b0000: BCD2 = 7'b1000000;
            4'b0001: BCD2 = 7'b1111001;
            4'b0010: BCD2 = 7'b0100100;
            4'b0011: BCD2 = 7'b0110000;
            4'b0100: BCD2 = 7'b0011001;
            4'b0101: BCD2 = 7'b0010010;
            4'b0110: BCD2 = 7'b0000010;
            4'b0111: BCD2 = 7'b1111000;
            4'b1000: BCD2 = 7'b0000000;
            4'b1001: BCD2 = 7'b0011000;
            4'b1010: BCD2 = 7'b0111111;
        endcase
        case(code[15:12])
            4'b0000: BCD3 = 7'b1000000;
            4'b0001: BCD3 = 7'b1111001;
            4'b0010: BCD3 = 7'b0100100;
            4'b0011: BCD3 = 7'b0110000;
            4'b0100: BCD3 = 7'b0011001;
            4'b0101: BCD3 = 7'b0010010;
            4'b0110: BCD3 = 7'b0000010;
            4'b0111: BCD3 = 7'b1111000;
            4'b1000: BCD3 = 7'b0000000;
            4'b1001: BCD3 = 7'b0011000;
            4'b1010: BCD3 = 7'b0111111;
        endcase
        case(code[19:16])
            4'b0000: BCD4 = 7'b1000000;
            4'b0001: BCD4 = 7'b1111001;
            4'b0010: BCD4 = 7'b0100100;
            4'b0011: BCD4 = 7'b0110000;
            4'b0100: BCD4 = 7'b0011001;
            4'b0101: BCD4 = 7'b0010010;
            4'b0110: BCD4 = 7'b0000010;
            4'b0111: BCD4 = 7'b1111000;
            4'b1000: BCD4 = 7'b0000000;
            4'b1001: BCD4 = 7'b0011000;
            4'b1010: BCD4 = 7'b0111111;
        endcase
        case(code[23:20])
            4'b0000: BCD5 = 7'b1000000;
            4'b0001: BCD5 = 7'b1111001;
            4'b0010: BCD5 = 7'b0100100;
            4'b0011: BCD5 = 7'b0110000;
            4'b0100: BCD5 = 7'b0011001;
            4'b0101: BCD5 = 7'b0010010;
            4'b0110: BCD5 = 7'b0000010;
            4'b0111: BCD5 = 7'b1111000;
            4'b1000: BCD5 = 7'b0000000;
            4'b1001: BCD5 = 7'b0011000;
            4'b1010: BCD5 = 7'b0111111;
        endcase
        case(code[27:24])
            4'b0000: BCD6 = 7'b1000000;
            4'b0001: BCD6 = 7'b1111001;
            4'b0010: BCD6 = 7'b0100100;
            4'b0011: BCD6 = 7'b0110000;
            4'b0100: BCD6 = 7'b0011001;
            4'b0101: BCD6 = 7'b0010010;
            4'b0110: BCD6 = 7'b0000010;
            4'b0111: BCD6 = 7'b1111000;
            4'b1000: BCD6 = 7'b0000000;
            4'b1001: BCD6 = 7'b0011000;
            4'b1010: BCD6 = 7'b0111111;
        endcase
end

endmodule